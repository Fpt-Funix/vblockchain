module io




fn test_create_blockchain() {

}
fn test_save_blockchain() {

	// create a new blockchain

	
	
}
fn test_save_then_load_blockchain() {

	
	
}
