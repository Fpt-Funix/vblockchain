module core

pub struct Transaction {
	hash string
	sender string
	recipient string
	amount int
	timestamp int
}
